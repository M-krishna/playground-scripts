module 4bitadder_tb;
    reg [3:0] in1;
    reg [3:0] in2;
    reg [3:0] out;
endmodule